`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/17/2017 02:21:06 PM
// Design Name: 
// Module Name: carry_pipe
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module d_ff ( a,b,c, clk, q,q1,q2);
   input a,b,c,clk;
   output q, q1,q2;
   wire clk;
   reg q, q1,q2;
     	 
   always @ (posedge clk)
   begin
    q <= a;
    q1<=b;
    q2 <= c;
 end

endmodule


module dff1 (s,cout,clk,q3,cout1);
   input s,clk,cout;
   output q3,cout1;
   wire clk;
   reg q3,cout1;
     	 
   always @ (posedge clk)
   begin
    q3 <= s;
    cout1 <= cout;
   
 end

endmodule


module carry_pipe(cout1,q3,a,b,cin,clk);
output [31:0]q3;
output cout1;
input [31:0]a,b;
input clk;
input cin;
wire [31:0]g,p,c,s;
wire cin1,cout;
wire [31:0]q,q1,q2,q3;

assign g=a&b;
assign p=a^b;

d_ff faa(a[0],b[0],cin,clk,q[0],q1[0],cin1);
assign c[0]=g[0]|(p[0]&cin);
d_ff f0(a[0],b[0],c[0],clk,q[0],q1[0],q2[0]);


assign c[1]=g[1]|(p[1]&(g[0]|(p[0]&cin)));
d_ff f1(a[1],b[1],c[1],clk,q[1],q1[1],q2[1]);

assign c[2]=g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))));
d_ff f2(a[2],b[2],c[2],clk,q[2],q1[2],q2[2]);

assign c[3]=g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))));
d_ff f3(a[3],b[3],c[3],clk,q[3],q1[3],q2[3]);

assign c[4]=g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))));
d_ff f4(a[4],b[4],c[4],clk,q[4],q1[4],q2[4]);

assign c[5]=g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))));
d_ff f5(a[5],b[5],c[5],clk,q[5],q1[5],q2[5]);

assign c[6]=g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))));
d_ff f6(a[6],b[6],c[6],clk,q[6],q1[6],q2[6]);

assign c[7]=g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))));
d_ff f7(a[7],b[7],c[7],clk,q[7],q1[7],q2[7]);

assign c[8]=g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))));
d_ff f8(a[8],b[8],c[8],clk,q[8],q1[8],q2[8]);

assign c[9]=g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))));
d_ff f9(a[9],b[9],c[9],clk,q[9],q1[9],q2[9]);

assign c[10]=g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))));
d_ff f10(a[10],b[10],c[10],clk,q[10],q1[10],q2[10]);

assign c[11]=g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))));
d_ff f11(a[11],b[11],c[11],clk,q[11],q1[11],q2[11]);

assign c[12]=g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))));
d_ff f12(a[12],b[12],c[12],clk,q[12],q1[12],q2[12]);

assign c[13]=g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))));
d_ff f13(a[13],b[13],c[13],clk,q[13],q1[13],q2[13]);

assign c[14]=g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))));
d_ff f14(a[14],b[14],c[14],clk,q[14],q1[14],q2[14]);

assign c[15]=g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))));
d_ff f15(a[15],b[15],c[15],clk,q[15],q1[15],q2[15]);

assign c[16]=g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))));
d_ff f16(a[16],b[16],c[16],clk,q[16],q1[16],q2[16]);

assign c[17]=g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))));
d_ff f17(a[17],b[17],c[17],clk,q[17],q1[17],q2[17]);

assign c[18]=g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))));
d_ff f18(a[18],b[18],c[18],clk,q[18],q1[18],q2[18]);

assign c[19]=g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))));
d_ff f19(a[19],b[19],c[19],clk,q[19],q1[19],q2[19]);

assign c[20]=g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))));
d_ff f20(a[20],b[20],c[20],clk,q[20],q1[20],q2[20]);

assign c[21]=g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))));
d_ff f21(a[21],b[21],c[21],clk,q[21],q1[21],q2[21]);

assign c[22]=g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))));
d_ff f22(a[22],b[22],c[22],clk,q[22],q1[22],q2[22]);

assign c[23]=g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))));
d_ff f23(a[23],b[23],c[23],clk,q[23],q1[23],q2[23]);

assign c[24]=g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f24(a[24],b[24],c[24],clk,q[24],q1[24],q2[24]);

assign c[25]=g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f25(a[25],b[25],c[25],clk,q[25],q1[25],q2[25]);

assign c[26]=g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p
[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f26(a[26],b[26],c[26],clk,q[26],q1[26],q2[26]);

assign c[27]=g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f27(a[27],b[27],c[27],clk,q[27],q1[27],q2[27]);

assign c[28]=g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f28(a[28],b[28],c[28],clk,q[28],q1[28],q2[28]);

assign c[29]=g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f29(a[29],b[29],c[29],clk,q[29],q1[29],q2[29]);

assign c[30]=g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f30(a[30],b[30],c[30],clk,q[30],q1[30],q2[30]);

assign c[31]=g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
d_ff f31(a[31],b[31],c[31],clk,q[31],q1[31],q2[31]);







assign s[0]=q[0]^q1[0]^cin1;
assign s[1]=q[1]^q1[1]^q2[0];
assign s[2]=q[2]^q1[2]^q2[1];
assign s[3]=q[3]^q1[3]^q2[2];
assign s[4]=q[4]^q1[4]^q2[3];
assign s[5]=q[5]^q1[5]^q2[4];
assign s[6]=q[6]^q1[6]^q2[5];
assign s[7]=q[7]^q1[7]^q2[6];
assign s[8]=q[8]^q1[8]^q2[7];
assign s[9]=q[9]^q1[9]^q2[8];
assign s[10]=q[10]^q1[10]^q2[9];
assign s[11]=q[11]^q1[11]^q2[10]; 
assign s[12]=q[12]^q1[12]^q2[11];
assign s[13]=q[13]^q1[13]^q2[12];
assign s[14]=q[14]^q1[14]^q2[13];
assign s[15]=q[15]^q1[15]^q2[14];
assign s[16]=q[16]^q1[16]^q2[15];
assign s[17]=q[17]^q1[17]^q2[16];
assign s[18]=q[18]^q1[18]^q2[17];
assign s[19]=q[19]^q1[19]^q2[18];
assign s[20]=q[20]^q1[20]^q2[19];
assign s[21]=q[21]^q1[21]^q2[20];
assign s[22]=q[22]^q1[22]^q2[21];
assign s[23]=q[23]^q1[23]^q2[22];
assign s[24]=q[24]^q1[24]^q2[23];
assign s[25]=q[25]^q1[25]^q2[24];
assign s[26]=q[26]^q1[26]^q2[25];
assign s[27]=q[27]^q1[27]^q2[26];
assign s[28]=q[28]^q1[28]^q2[27];
assign s[29]=q[29]^q1[29]^q2[28];
assign s[30]=q[30]^q1[30]^q2[29];
assign s[31]=q[31]^q1[31]^q2[30];
assign cout=q2[31];

dff1 ob(s[0],cout,clk,q3[0],cout1);
dff1 ob1(s[1],cout,clk,q3[1],cout1);
dff1 ob2(s[2],cout,clk,q3[2],cout1);
dff1 ob3(s[3],cout,clk,q3[3],cout1);
dff1 ob111(s[4],cout,clk,q3[4],cout1);
dff1 ob4(s[5],cout,clk,q3[5],cout1);
dff1 ob5(s[6],cout,clk,q3[6],cout1);
dff1 ob6(s[7],cout,clk,q3[7],cout1);
dff1 ob7(s[8],cout,clk,q3[8],cout1);
dff1 ob8(s[9],cout,clk,q3[9],cout1);
dff1 ob9(s[10],cout,clk,q3[10],cout1);
dff1 ob10(s[11],cout,clk,q3[11],cout1);
dff1 ob11(s[12],cout,clk,q3[12],cout1);
dff1 ob12(s[13],cout,clk,q3[13],cout1);
dff1 ob13(s[14],cout,clk,q3[14],cout1);
dff1 ob14(s[15],cout,clk,q3[15],cout1);
dff1 ob15(s[16],cout,clk,q3[16],cout1);
dff1 ob16(s[17],cout,clk,q3[17],cout1);
dff1 ob17(s[18],cout,clk,q3[18],cout1);
dff1 ob18(s[19],cout,clk,q3[19],cout1);
dff1 ob19(s[20],cout,clk,q3[20],cout1);
dff1 ob20(s[21],cout,clk,q3[21],cout1);
dff1 ob21(s[22],cout,clk,q3[22],cout1);
dff1 ob22(s[23],cout,clk,q3[23],cout1);
dff1 ob23(s[24],cout,clk,q3[24],cout1);
dff1 ob24(s[25],cout,clk,q3[25],cout1);
dff1 ob25(s[26],cout,clk,q3[26],cout1);
dff1 ob26(s[27],cout,clk,q3[27],cout1);
dff1 ob27(s[28],cout,clk,q3[28],cout1);
dff1 ob28(s[29],cout,clk,q3[29],cout1);
dff1 ob29(s[30],cout,clk,q3[30],cout1);
dff1 ob30(s[31],cout,clk,q3[31],cout1);





endmodule





