module main(sa,sb,ea,eb,ma,mb,ma_out,signbit,exponent,clk);
input [22:0]ma,mb;
input sa,sb;
input [7:0]ea,eb;

output reg [23:0]ma_out;
 reg result;
output signbit;
input clk;
output [7:0]exponent;
wire [31:0]ma1,mb1;
wire [63:0]R;
wire [8:0]exp1;
wire [8:0]ea1,eb1,exp;
wire [8:0]subt;
wire cout,cout1;
assign ma1[22:0]=ma[22:0];
assign ma1[23]=1'b1;
assign ma1[31:24]=8'b0;

assign mb1[22:0]=mb[22:0];
assign mb1[23]=1'b1;
assign mb1[31:24]=8'b0;

wallacetreemult maaaa(ma1,mb1,R,carry,clk);

always@(*)
begin
if(R[46]==1'b1)
begin
	ma_out[23:0]<=R[47:23];
	result<=R[47];
	
end
else if(R[47]==1'b1)
begin
	ma_out[23:0]<=R[48:24];
	//ma_out[23]<=R[47];
	
end
end

assign signbit=sa^sb;

assign ea1[7:0]=ea[7:0];
assign ea1[8]=1'b0;

assign eb1[7:0]=eb[7:0];
assign eb1[8]=1'b0;

cla9 chjkl(cout,exp,ea1,eb1,0);


assign subt=9'd127;

cla9 cabg(cout1,exp1,exp,~subt,1);

assign exponent[7:0]=exp1[7:0];

endmodule

module cla9(cout,s,a,b,cin);

input [8:0]a,b;
input cin;

output [8:0]s;
output cout;
wire [8:0]g,p,c;
assign g=a&b;
assign p=a^b;
assign c[0]=g[0]|(p[0]&cin);
assign c[1]=g[1]|(p[1]&(g[0]|(p[0]&cin)));
assign c[2]=g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))));
assign c[3]=g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))));
assign c[4]=g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))));

assign c[5]=g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))));

assign c[6]=g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))));

assign c[7]=g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))));

assign c[8]=g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))));

assign cout=c[8];

assign s[0]=p[0]^cin;
assign s[1]=p[1]^c[0];
assign s[2]=p[2]^c[1];
assign s[3]=p[3]^c[2];
assign s[4]=p[4]^c[3];
assign s[5]=p[5]^c[4];
assign s[6]=p[6]^c[5];
assign s[7]=p[7]^c[6];
assign s[8]=p[8]^c[7];


endmodule

//`include "csa.v"
//`include "cla32.v"
//`include "ff.v"
module wallacetreemult(A,B,R,carry,clk);
input [31:0]A,B;
input clk;
wire [63:0]U[63:0];
wire [63:0]V[63:0];
output [63:0]R;
output carry;
wire [63:0]P[63:0];
wire [63:0]q[63:0];
wire [63:0]q1[63:0];
wire [63:0]p1[63:0];


assign P[0]=B[0]?{32'b000,A}:64'h0000;
assign P[1]=B[1]?{32'b000,A}<<1:64'h0000;
assign P[2]=B[2]?{32'b000,A}<<2:64'h0000;
assign P[3]=B[3]?{32'b000,A}<<3:64'h0000;
assign P[4]=B[4]?{32'b000,A}<<4:64'h0000;
assign P[5]=B[5]?{32'b000,A}<<5:64'h0000;
assign P[6]=B[6]?{32'b000,A}<<6:64'h0000;
assign P[7]=B[7]?{32'b000,A}<<7:64'h0000;

assign P[8]=B[8]?{32'b000,A}<<8:64'h0000;
assign P[9]=B[9]?{32'b000,A}<<9:64'h0000;
assign P[10]=B[10]?{32'b000,A}<<10:64'h0000;
assign P[11]=B[11]?{32'b000,A}<<11:64'h0000;
assign P[12]=B[12]?{32'b000,A}<<12:64'h0000;
assign P[13]=B[13]?{32'b000,A}<<13:64'h0000;
assign P[14]=B[14]?{32'b000,A}<<14:64'h0000;
assign P[15]=B[15]?{32'b000,A}<<15:64'h0000;

assign P[16]=B[16]?{32'b000,A}<<16:64'h0000;
assign P[17]=B[17]?{32'b000,A}<<17:64'h0000;
assign P[18]=B[18]?{32'b000,A}<<18:64'h0000;
assign P[19]=B[19]?{32'b000,A}<<19:64'h0000;
assign P[20]=B[20]?{32'b000,A}<<20:64'h0000;
assign P[21]=B[21]?{32'b000,A}<<21:64'h0000;
assign P[22]=B[22]?{32'b000,A}<<22:64'h0000;
assign P[23]=B[23]?{32'b000,A}<<23:64'h0000;

assign P[24]=B[24]?{32'b000,A}<<24:64'h0000;
assign P[25]=B[25]?{32'b000,A}<<25:64'h0000;
assign P[26]=B[26]?{32'b000,A}<<26:64'h0000;
assign P[27]=B[27]?{32'b000,A}<<27:64'h0000;
assign P[28]=B[28]?{32'b000,A}<<28:64'h0000;
assign P[29]=B[29]?{32'b000,A}<<29:64'h0000;
assign P[30]=B[30]?{32'b000,A}<<30:64'h0000;
assign P[31]=B[31]?{32'b000,A}<<31:64'h0000;

//1ssst
csaveadder c1(P[0],P[1],P[2],U[0],V[0]);
d_ff f0 ( U[0],V[0], clk, q[0],q1[0]);

csaveadder c2(P[3],P[4],P[5],U[1],V[1]);
d_ff f1 ( U[1],V[1], clk, q[1],q1[1]);

csaveadder c3(P[6],P[7],P[8],U[2],V[2]);
d_ff f2 ( U[2],V[2], clk, q[2],q1[2]);

csaveadder c4(P[9],P[10],P[11],U[3],V[3]);
d_ff f3 ( U[3],V[3], clk, q[3],q1[3]);

csaveadder c5(P[12],P[13],P[14],U[4],V[4]);
d_ff f4 ( U[4],V[4], clk, q[4],q1[4]);

csaveadder c6(P[15],P[16],P[17],U[5],V[5]);
d_ff f5 ( U[5],V[5], clk, q[5],q1[5]);

csaveadder c7(P[18],P[19],P[20],U[6],V[6]);
d_ff f6 ( U[6],V[6], clk, q[6],q1[6]);

csaveadder c8(P[21],P[22],P[23],U[7],V[7]);
d_ff f7 ( U[7],V[7], clk, q[7],q1[7]);

csaveadder c9(P[24],P[25],P[26],U[8],V[8]);
d_ff f8 ( U[8],V[8], clk, q[8],q1[8]);

csaveadder c10(P[27],P[28],P[29],U[9],V[9]);
d_ff f9 ( U[9],V[9], clk, q[9],q1[9]);

d_ff f10( P[30],P[31],clk,p1[1],p1[2]);
//

//2ndd
csaveadder c11(q[0],q1[0],q[1],U[10],V[10]);
d_ff f11 ( U[10],V[10], clk, q[10],q1[10]);
 
csaveadder c12(q1[1],q[2],q1[2],U[11],V[11]);
d_ff f12 ( U[11],V[11], clk, q[11],q1[11]);

csaveadder c13(q[3],q1[3],q[4],U[12],V[12]);
d_ff f13 ( U[12],V[12], clk, q[12],q1[12]);

csaveadder c14(q1[4],q[5],q1[5],U[13],V[13]);
d_ff f14 ( U[13],V[13], clk, q[13],q1[13]);

csaveadder c15(q[6],q1[6],q[7],U[14],V[14]);
d_ff f15 ( U[14],V[14], clk, q[14],q1[14]);

csaveadder c16(q1[7],q[8],q1[8],U[15],V[15]);
d_ff f16 ( U[15],V[15], clk, q[15],q1[15]);

csaveadder c17(q[9],q1[9],p1[1],U[16],V[16]);
d_ff f17 ( U[16],V[16], clk, q[16],q1[16]);

d_ff f18 ( p1[2],p1[2],clk,p1[3],p1[4]);//p1[3]=p1[4]
//


//3rdd
csaveadder c18(q[10],q1[10],q[11],U[17],V[17]);
d_ff f19 ( U[17],V[17], clk, q[17],q1[17]);

csaveadder c19(q1[11],q[12],q1[12],U[18],V[18]);
d_ff f20 ( U[18],V[18], clk, q[18],q1[18]);

csaveadder c20(q[13],q1[13],q[14],U[19],V[19]);
d_ff f21 ( U[19],V[19], clk, q[19],q1[19]);

csaveadder c21(q1[14],q[15],q1[15],U[20],V[20]);
d_ff f22 ( U[20],V[20], clk, q[20],q1[20]);

csaveadder c22(q[16],q1[16],p1[4],U[21],V[21]);//p1[3]=p[31]
d_ff f23 ( U[21],V[21], clk, q[21],q1[21]);

d_ff f24 ( V[21],V[21], clk, p1[5],p1[6]);
//


//4th
csaveadder c23(q[17],q1[17],q[18],U[22],V[22]);
d_ff f25 ( U[22],V[22], clk, q[22],q1[22]);

csaveadder c24(q1[18],q[19],q1[19],U[23],V[23]);
d_ff f26 ( U[23],V[23], clk, q[23],q1[23]);

csaveadder c25(q[20],q1[20],q[21],U[24],V[24]);
d_ff f27 ( U[24],V[24], clk, q[24],q1[24]);

d_ff f28 ( p1[5],p1[6], clk, p1[7],p1[8]);
//


//5thhh

csaveadder c26(q[22],q1[22],q[23],U[25],V[25]);
d_ff f29 ( U[25],V[25], clk, q[25],q1[25]);

csaveadder c27(q1[23],q[24],q1[24],U[26],V[26]);
d_ff f30 ( U[26],V[26], clk, q[26],q1[26]);

d_ff f31 ( p1[7],p1[8], clk, p1[9],p1[10]);
//


//6thh
csaveadder c28(q[25],q1[25],q[26],U[27],V[27]);
d_ff f32 ( U[27],V[27], clk, q[27],q1[27]);

d_ff f33 ( p1[9],p1[10], clk, p1[11],p1[12]);
//


//7thh
csaveadder c29(q1[26],q[27],q1[27],U[28],V[28]);
d_ff f34 ( U[28],V[28], clk, q[28],q1[28]);

d_ff f35 ( p1[11],p1[12], clk, p1[13],p1[14]);

//


//8thh
csaveadder c30(q[28],q1[28],p1[13],U[29],V[29]);
d_ff f36 ( U[29],V[29], clk, q[29],q1[29]);

//
//rca_64bit q0(q[29],q1[29],0,R,carry);
cla32 c000(carry,R,q[29],q1[29],0);
//cla32(cout,s,a,b,cin);
endmodule


module fulladder(a,b,cin,s,cout);

input a,b,cin;
output s,cout;

assign s=a^b^cin;
assign cout=(a&b)|(b&cin)|(a&cin);

endmodule


//`include "fa.v"
module csaveadder(X,Y,Z,U,V);
input [63:0]X;
input [63:0]Y;
input [63:0]Z;
output [63:0]U;
output [63:0]V;
wire temp;

assign V[0]=0;

fulladder fa0(X[0],Y[0],Z[0],U[0],V[1]);
fulladder fa1(X[1],Y[1],Z[1],U[1],V[2]);
fulladder fa2(X[2],Y[2],Z[2],U[2],V[3]);
fulladder fa3(X[3],Y[3],Z[3],U[3],V[4]);
fulladder fa4(X[4],Y[4],Z[4],U[4],V[5]);
fulladder fa5(X[5],Y[5],Z[5],U[5],V[6]);
fulladder fa6(X[6],Y[6],Z[6],U[6],V[7]);
fulladder fa7(X[7],Y[7],Z[7],U[7],V[8]);
fulladder fa8(X[8],Y[8],Z[8],U[8],V[9]);
fulladder fa9(X[9],Y[9],Z[9],U[9],V[10]);
fulladder fa10(X[10],Y[10],Z[10],U[10],V[11]);
fulladder fa11(X[11],Y[11],Z[11],U[11],V[12]);
fulladder fa12(X[12],Y[12],Z[12],U[12],V[13]);
fulladder fa13(X[13],Y[13],Z[13],U[13],V[14]);
fulladder fa14(X[14],Y[14],Z[14],U[14],V[15]);
fulladder fa15(X[15],Y[15],Z[15],U[15],V[16]);
fulladder fa16(X[16],Y[16],Z[16],U[16],V[17]);
fulladder fa17(X[17],Y[17],Z[17],U[17],V[18]);
fulladder fa18(X[18],Y[18],Z[18],U[18],V[19]);
fulladder fa19(X[19],Y[19],Z[19],U[19],V[20]);
fulladder fa20(X[20],Y[20],Z[20],U[20],V[21]);
fulladder fa21(X[21],Y[21],Z[21],U[21],V[22]);
fulladder fa22(X[22],Y[22],Z[22],U[22],V[23]);
fulladder fa23(X[23],Y[23],Z[23],U[23],V[24]);
fulladder fa24(X[24],Y[24],Z[24],U[24],V[25]);
fulladder fa25(X[25],Y[25],Z[25],U[25],V[26]);
fulladder fa26(X[26],Y[26],Z[26],U[26],V[27]);
fulladder fa27(X[27],Y[27],Z[27],U[27],V[28]);
fulladder fa28(X[28],Y[28],Z[28],U[28],V[29]);
fulladder fa29(X[29],Y[29],Z[29],U[29],V[30]);
fulladder fa30(X[30],Y[30],Z[30],U[30],V[31]);
fulladder fa31(X[31],Y[31],Z[31],U[31],V[32]);
fulladder fa32(X[32],Y[32],Z[32],U[32],V[33]);
fulladder fa33(X[33],Y[33],Z[33],U[33],V[34]);
fulladder fa34(X[34],Y[34],Z[34],U[34],V[35]);
fulladder fa35(X[35],Y[35],Z[35],U[35],V[36]);
fulladder fa36(X[36],Y[36],Z[36],U[36],V[37]);
fulladder fa37(X[37],Y[37],Z[37],U[37],V[38]);
fulladder fa38(X[38],Y[38],Z[38],U[38],V[39]);
fulladder fa39(X[39],Y[39],Z[39],U[39],V[40]);
fulladder fa40(X[40],Y[40],Z[40],U[40],V[41]);
fulladder fa41(X[41],Y[41],Z[41],U[41],V[42]);
fulladder fa42(X[42],Y[42],Z[42],U[42],V[43]);
fulladder fa43(X[43],Y[43],Z[43],U[43],V[44]);
fulladder fa44(X[44],Y[44],Z[44],U[44],V[45]);
fulladder fa45(X[45],Y[45],Z[45],U[45],V[46]);
fulladder fa46(X[46],Y[46],Z[46],U[46],V[47]);
fulladder fa47(X[47],Y[47],Z[47],U[47],V[48]);
fulladder fa48(X[48],Y[48],Z[48],U[48],V[49]);
fulladder fa49(X[49],Y[49],Z[49],U[49],V[50]);
fulladder fa50(X[50],Y[50],Z[50],U[50],V[51]);
fulladder fa51(X[51],Y[51],Z[51],U[51],V[52]);
fulladder fa52(X[52],Y[52],Z[52],U[52],V[53]);
fulladder fa53(X[53],Y[53],Z[53],U[53],V[54]);
fulladder fa54(X[54],Y[54],Z[54],U[54],V[55]);
fulladder fa55(X[55],Y[55],Z[55],U[55],V[56]);
fulladder fa56(X[56],Y[56],Z[56],U[56],V[57]);
fulladder fa57(X[57],Y[57],Z[57],U[57],V[58]);
fulladder fa58(X[58],Y[58],Z[58],U[58],V[59]);
fulladder fa59(X[59],Y[59],Z[59],U[59],V[60]);
fulladder fa60(X[60],Y[60],Z[60],U[60],V[61]);
fulladder fa61(X[61],Y[61],Z[61],U[61],V[62]);
fulladder fa62(X[62],Y[62],Z[62],U[62],V[63]);
fulladder fa63(X[63],Y[63],Z[63],U[63],temp);

endmodule

module d_ff ( a,b, clk, q,q1);
   input [63:0]a;
   input [63:0]b;
   //input [63:0]c;
   input clk;
   output [63:0]q;
   output  [63:0]q1;	
  // output [63:0]q63;
   wire clk;
   reg [63:0]q;
   reg  [63:0]q1;
   //reg [63:0]q63;
   always @ (posedge clk)
   begin
    q <= a;
    q1 <=b;
    //q63 <= c;
 end

endmodule

//`include "ff.v"
//`include "dff1.v"
module cla32(cout,s,a,b,cin);
output [63:0]s;
output cout;
input [63:0]a,b;
//input clk;
input cin;
wire [63:0]g,p,c,s;
//wire cin1,cout;
//wire [31:0]q,b,c,q3;

assign g=a&b;
assign p=a^b;

//d_ff faa(a[0],b[0],cin,clk,q[0],b[0],cin1);
assign c[0]=g[0]|(p[0]&cin);
//d_ff f0(a[0],b[0],c[0],clk,q[0],b[0],c[0]);


assign c[1]=g[1]|(p[1]&(g[0]|(p[0]&cin)));
//d_ff f1(a[1],b[1],c[1],clk,q[1],b[1],c[1]);

assign c[2]=g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))));
//d_ff f2(a[2],b[2],c[2],clk,q[2],b[2],c[2]);

assign c[3]=g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))));
//d_ff f3(a[3],b[3],c[3],clk,q[3],b[3],c[3]);

assign c[4]=g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))));
//d_ff f4(a[4],b[4],c[4],clk,q[4],b[4],c[4]);

assign c[5]=g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))));
//d_ff f5(a[5],b[5],c[5],clk,q[5],b[5],c[5]);

assign c[6]=g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))));
//d_ff f6(a[6],b[6],c[6],clk,q[6],b[6],c[6]);

assign c[7]=g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))));
//d_ff f7(a[7],b[7],c[7],clk,q[7],b[7],c[7]);

assign c[8]=g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))));
//d_ff f8(a[8],b[8],c[8],clk,q[8],b[8],c[8]);

assign c[9]=g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))));
//d_ff f9(a[9],b[9],c[9],clk,q[9],b[9],c[9]);

assign c[10]=g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))));
//d_ff f10(a[10],b[10],c[10],clk,q[10],b[10],c[10]);

assign c[11]=g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))));
//d_ff f11(a[11],b[11],c[11],clk,q[11],b[11],c[11]);

assign c[12]=g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))));
//d_ff f12(a[12],b[12],c[12],clk,q[12],b[12],c[12]);

assign c[13]=g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))));
//d_ff f13(a[13],b[13],c[13],clk,q[13],b[13],c[13]);

assign c[14]=g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))));
//d_ff f14(a[14],b[14],c[14],clk,q[14],b[14],c[14]);

assign c[15]=g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))));
//d_ff f15(a[15],b[15],c[15],clk,q[15],b[15],c[15]);

assign c[16]=g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))));
//d_ff f16(a[16],b[16],c[16],clk,q[16],b[16],c[16]);

assign c[17]=g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))));
//d_ff f17(a[17],b[17],c[17],clk,q[17],b[17],c[17]);

assign c[18]=g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))));
//d_ff f18(a[18],b[18],c[18],clk,q[18],b[18],c[18]);

assign c[19]=g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))));
//d_ff f19(a[19],b[19],c[19],clk,q[19],b[19],c[19]);

assign c[20]=g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))));
//d_ff f20(a[20],b[20],c[20],clk,q[20],b[20],c[20]);

assign c[21]=g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))));
//d_ff f21(a[21],b[21],c[21],clk,q[21],b[21],c[21]);

assign c[22]=g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))));
//d_ff f22(a[22],b[22],c[22],clk,q[22],b[22],c[22]);

assign c[23]=g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f23(a[23],b[23],c[23],clk,q[23],b[23],c[23]);

assign c[24]=g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f24(a[24],b[24],c[24],clk,q[24],b[24],c[24]);

assign c[25]=g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f25(a[25],b[25],c[25],clk,q[25],b[25],c[25]);

assign c[26]=g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p
[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f26(a[26],b[26],c[26],clk,q[26],b[26],c[26]);

assign c[27]=g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f27(a[27],b[27],c[27],clk,q[27],b[27],c[27]);

assign c[28]=g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f28(a[28],b[28],c[28],clk,q[28],b[28],c[28]);

assign c[29]=g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f29(a[29],b[29],c[29],clk,q[29],b[29],c[29]);

assign c[30]=g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f30(a[30],b[30],c[30],clk,q[30],b[30],c[30]);

assign c[31]=g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
//d_ff f31(a[31],b[31],c[31],clk,q[31],b[31],c[31]);

assign c[32]=g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[33]=g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[34]=g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[35]=g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[36]=g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[37]=g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[38]=g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[39]=g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[40]=g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[41]=g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[42]=g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[43]=g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[44]=g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[45]=g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[46]=g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[47]=g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[48]=g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[49]=g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[50]=g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[51]=g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[52]=g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[53]=g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[54]=g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[55]=g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


assign c[56]=g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[57]=g[57]|(p[57]&(g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[58]=g[58]|(p[58]&(g[57]|(p[57]&(g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[59]=g[59]|(p[59]&(g[58]|(p[58]&(g[57]|(p[57]&(g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[60]=g[60]|(p[60]&(g[59]|(p[59]&(g[58]|(p[58]&(g[57]|(p[57]&(g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[61]=g[61]|(p[61]&(g[60]|(p[60]&(g[59]|(p[59]&(g[58]|(p[58]&(g[57]|(p[57]&(g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[62]=g[62]|(p[62]&(g[61]|(p[61]&(g[60]|(p[60]&(g[59]|(p[59]&(g[58]|(p[58]&(g[57]|(p[57]&(g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[63]=g[63]|(p[63]&(g[62]|(p[62]&(g[61]|(p[61]&(g[60]|(p[60]&(g[59]|(p[59]&(g[58]|(p[58]&(g[57]|(p[57]&(g[56]|(p[56]&(g[55]|(p[55]&(g[54]|(p[54]&(g[53]|(p[53]&(g[52]|(p[51]&(g[51]|(p[51]&(g[50]|(p[50]&(g[49]|(p[49]&(g[48]|(p[48]&(g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(g[20]&(g[19]|(p[19]&g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));




assign s[0]=a[0]^b[0]^cin;
assign s[1]=a[1]^b[1]^c[0];
assign s[2]=a[2]^b[2]^c[1];
assign s[3]=a[3]^b[3]^c[2];
assign s[4]=a[4]^b[4]^c[3];
assign s[5]=a[5]^b[5]^c[4];
assign s[6]=a[6]^b[6]^c[5];
assign s[7]=a[7]^b[7]^c[6];
assign s[8]=a[8]^b[8]^c[7];
assign s[9]=a[9]^b[9]^c[8];
assign s[10]=a[10]^b[10]^c[9];
assign s[11]=a[11]^b[11]^c[10]; 
assign s[12]=a[12]^b[12]^c[11];
assign s[13]=a[13]^b[13]^c[12];
assign s[14]=a[14]^b[14]^c[13];
assign s[15]=a[15]^b[15]^c[14];
assign s[16]=a[16]^b[16]^c[15];
assign s[17]=a[17]^b[17]^c[16];
assign s[18]=a[18]^b[18]^c[17];
assign s[19]=a[19]^b[19]^c[18];
assign s[20]=a[20]^b[20]^c[19];
assign s[21]=a[21]^b[21]^c[20];
assign s[22]=a[22]^b[22]^c[21];
assign s[23]=a[23]^b[23]^c[22];
assign s[24]=a[24]^b[24]^c[23];
assign s[25]=a[25]^b[25]^c[24];
assign s[26]=a[26]^b[26]^c[25];
assign s[27]=a[27]^b[27]^c[26];
assign s[28]=a[28]^b[28]^c[27];
assign s[29]=a[29]^b[29]^c[28];
assign s[30]=a[30]^b[30]^c[29];
assign s[31]=a[31]^b[31]^c[30];
assign s[32]=a[32]^b[32]^c[31];
assign s[33]=a[33]^b[33]^c[32];
assign s[34]=a[34]^b[34]^c[33];
assign s[35]=a[35]^b[35]^c[34];
assign s[36]=a[36]^b[36]^c[35];
assign s[37]=a[37]^b[37]^c[36];
assign s[38]=a[38]^b[38]^c[37];
assign s[39]=a[39]^b[39]^c[38];
assign s[40]=a[40]^b[40]^c[39];
assign s[41]=a[41]^b[41]^c[40];
assign s[42]=a[42]^b[42]^c[41];
assign s[43]=a[43]^b[43]^c[42];
assign s[44]=a[44]^b[44]^c[43];
assign s[45]=a[45]^b[45]^c[44];
assign s[46]=a[46]^b[46]^c[45];
assign s[47]=a[47]^b[47]^c[46];
assign s[48]=a[48]^b[48]^c[47];
assign s[49]=a[49]^b[49]^c[48];
assign s[50]=a[50]^b[50]^c[49];
assign s[51]=a[51]^b[51]^c[50];
assign s[52]=a[52]^b[52]^c[51];
assign s[53]=a[53]^b[53]^c[52];
assign s[54]=a[54]^b[54]^c[53];
assign s[55]=a[55]^b[55]^c[54];
assign s[56]=a[56]^b[56]^c[55];
assign s[57]=a[57]^b[57]^c[56];
assign s[58]=a[58]^b[58]^c[57];
assign s[59]=a[59]^b[59]^c[58];
assign s[60]=a[60]^b[60]^c[59];
assign s[61]=a[61]^b[61]^c[60];
assign s[62]=a[62]^b[62]^c[61];
assign s[63]=a[63]^b[63]^c[62];

assign cout=c[63];





endmodule

